`timescale 1ns /1ps
///////////////////////////////////////////////////////////////////
// Authored by David J. Marion aka FPGA Dude
// Created on 4/13/2022
//
// Description: ROM containing 8x16 ascii characters for clock
// and calendar on VGA
///////////////////////////////////////////////////////////////////

module clock_digit_rom(
   input clk, 
   input wire [10:0] addr,
   output reg [7:0] data
   );
    
   (* rom_style = "block" *)   

   reg [10:0] addr_reg;
   
   always @(posedge clk)
      addr_reg <= addr;
      
   always @*
      case(addr_reg)
        // code x2e (.)
         11'h2e0: data = 8'b00000000;   //
         11'h2e1: data = 8'b00000000;   //
         11'h2e2: data = 8'b00000000;   //
         11'h2e3: data = 8'b00000000;   //
         11'h2e4: data = 8'b00000000;   //
         11'h2e5: data = 8'b00000000;   //
         11'h2e6: data = 8'b00000000;   //
         11'h2e7: data = 8'b00000000;   //
         11'h2e8: data = 8'b00000000;   //
         11'h2e9: data = 8'b00000000;   //
         11'h2ea: data = 8'b00011000;   //   **
         11'h2eb: data = 8'b00011000;   //   **
         11'h2ec: data = 8'b00000000;   //
         11'h2ed: data = 8'b00000000;   //
         11'h2ee: data = 8'b00000000;   //
         11'h2ef: data = 8'b00000000;   //
         // code x30 (0)
         11'h300: data = 8'b00000000;   //
         11'h301: data = 8'b00000000;   //
         11'h302: data = 8'b00111000;   //  ***  
         11'h303: data = 8'b01101100;   // ** **
         11'h304: data = 8'b11000110;   //**   **
         11'h305: data = 8'b11000110;   //**   **
         11'h306: data = 8'b11000110;   //**   **
         11'h307: data = 8'b11000110;   //**   **
         11'h308: data = 8'b11000110;   //**   **
         11'h309: data = 8'b11000110;   //**   **
         11'h30a: data = 8'b01101100;   // ** **
         11'h30b: data = 8'b00111000;   //  ***
         11'h30c: data = 8'b00000000;   //
         11'h30d: data = 8'b00000000;   //
         11'h30e: data = 8'b00000000;   //
         11'h30f: data = 8'b00000000;   //
         // code x31 (1)
         11'h310: data = 8'b00000000;   //
         11'h311: data = 8'b00000000;   //
         11'h312: data = 8'b00011000;   //   **  
         11'h313: data = 8'b00111000;   //  ***
         11'h314: data = 8'b01111000;   // ****
         11'h315: data = 8'b00011000;   //   **
         11'h316: data = 8'b00011000;   //   **
         11'h317: data = 8'b00011000;   //   **
         11'h318: data = 8'b00011000;   //   **
         11'h319: data = 8'b00011000;   //   **
         11'h31a: data = 8'b01111110;   // ******
         11'h31b: data = 8'b01111110;   // ******
         11'h31c: data = 8'b00000000;   //
         11'h31d: data = 8'b00000000;   //
         11'h31e: data = 8'b00000000;   //
         11'h31f: data = 8'b00000000;   //
         // code x32 (2)
         11'h320: data = 8'b00000000;   //
         11'h321: data = 8'b00000000;   //
         11'h322: data = 8'b11111110;   //*******  
         11'h323: data = 8'b11111110;   //*******
         11'h324: data = 8'b00000110;   //     **
         11'h325: data = 8'b00000110;   //     **
         11'h326: data = 8'b11111110;   //*******
         11'h327: data = 8'b11111110;   //*******
         11'h328: data = 8'b11000000;   //**
         11'h329: data = 8'b11000000;   //**
         11'h32a: data = 8'b11111110;   //*******
         11'h32b: data = 8'b11111110;   //*******
         11'h32c: data = 8'b00000000;   //
         11'h32d: data = 8'b00000000;   //
         11'h32e: data = 8'b00000000;   //
         11'h32f: data = 8'b00000000;   //
         // code x33 (3)
         11'h330: data = 8'b00000000;   //
         11'h331: data = 8'b00000000;   //
         11'h332: data = 8'b11111110;   //*******  
         11'h333: data = 8'b11111110;   //*******
         11'h334: data = 8'b00000110;   //     **
         11'h335: data = 8'b00000110;   //     **
         11'h336: data = 8'b00111110;   //  *****
         11'h337: data = 8'b00111110;   //  *****
         11'h338: data = 8'b00000110;   //     **
         11'h339: data = 8'b00000110;   //     **
         11'h33a: data = 8'b11111110;   //*******
         11'h33b: data = 8'b11111110;   //*******
         11'h33c: data = 8'b00000000;   //
         11'h33d: data = 8'b00000000;   //
         11'h33e: data = 8'b00000000;   //
         11'h33f: data = 8'b00000000;   //
         // code x34 (4)
         11'h340: data = 8'b00000000;   //
         11'h341: data = 8'b00000000;   //
         11'h342: data = 8'b11000110;   //**   **  
         11'h343: data = 8'b11000110;   //**   **
         11'h344: data = 8'b11000110;   //**   **
         11'h345: data = 8'b11000110;   //**   **
         11'h346: data = 8'b11111110;   //*******
         11'h347: data = 8'b11111110;   //*******
         11'h348: data = 8'b00000110;   //     **
         11'h349: data = 8'b00000110;   //     **
         11'h34a: data = 8'b00000110;   //     **
         11'h34b: data = 8'b00000110;   //     **
         11'h34c: data = 8'b00000000;   //
         11'h34d: data = 8'b00000000;   //
         11'h34e: data = 8'b00000000;   //
         11'h34f: data = 8'b00000000;   //
         // code x35 (5)
         11'h350: data = 8'b00000000;   //
         11'h351: data = 8'b00000000;   //
         11'h352: data = 8'b11111110;   //*******  
         11'h353: data = 8'b11111110;   //*******
         11'h354: data = 8'b11000000;   //**
         11'h355: data = 8'b11000000;   //**
         11'h356: data = 8'b11111110;   //*******
         11'h357: data = 8'b11111110;   //*******
         11'h358: data = 8'b00000110;   //     **
         11'h359: data = 8'b00000110;   //     **
         11'h35a: data = 8'b11111110;   //*******
         11'h35b: data = 8'b11111110;   //*******
         11'h35c: data = 8'b00000000;   //
         11'h35d: data = 8'b00000000;   //
         11'h35e: data = 8'b00000000;   //
         11'h35f: data = 8'b00000000;   //
         // code x36 (6)
         11'h360: data = 8'b00000000;   //
         11'h361: data = 8'b00000000;   //
         11'h362: data = 8'b11111110;   //*******  
         11'h363: data = 8'b11111110;   //*******
         11'h364: data = 8'b11000000;   //**
         11'h365: data = 8'b11000000;   //**
         11'h366: data = 8'b11111110;   //*******
         11'h367: data = 8'b11111110;   //*******
         11'h368: data = 8'b11000110;   //**   **
         11'h369: data = 8'b11000110;   //**   **
         11'h36a: data = 8'b11111110;   //*******
         11'h36b: data = 8'b11111110;   //*******
         11'h36c: data = 8'b00000000;   //
         11'h36d: data = 8'b00000000;   //
         11'h36e: data = 8'b00000000;   //
         11'h36f: data = 8'b00000000;   //
         // code x37 (7)
         11'h370: data = 8'b00000000;   //
         11'h371: data = 8'b00000000;   //
         11'h372: data = 8'b11111110;   //*******  
         11'h373: data = 8'b11111110;   //*******
         11'h374: data = 8'b00000110;   //     **
         11'h375: data = 8'b00000110;   //     **
         11'h376: data = 8'b00000110;   //     **
         11'h377: data = 8'b00000110;   //     **
         11'h378: data = 8'b00000110;   //     **
         11'h379: data = 8'b00000110;   //     **
         11'h37a: data = 8'b00000110;   //     **
         11'h37b: data = 8'b00000110;   //     **
         11'h37c: data = 8'b00000000;   //
         11'h37d: data = 8'b00000000;   //
         11'h37e: data = 8'b00000000;   //
         11'h37f: data = 8'b00000000;   //
         // code x38 (8)
         11'h380: data = 8'b00000000;   //
         11'h381: data = 8'b00000000;   //
         11'h382: data = 8'b11111110;   //*******  
         11'h383: data = 8'b11111110;   //*******
         11'h384: data = 8'b11000110;   //**   **
         11'h385: data = 8'b11000110;   //**   **
         11'h386: data = 8'b11111110;   //*******
         11'h387: data = 8'b11111110;   //*******
         11'h388: data = 8'b11000110;   //**   **
         11'h389: data = 8'b11000110;   //**   **
         11'h38a: data = 8'b11111110;   //*******
         11'h38b: data = 8'b11111110;   //*******
         11'h38c: data = 8'b00000000;   //
         11'h38d: data = 8'b00000000;   //
         11'h38e: data = 8'b00000000;   //
         11'h38f: data = 8'b00000000;   //
         // code x39 (9)
         11'h390: data = 8'b00000000;   //
         11'h391: data = 8'b00000000;   //
         11'h392: data = 8'b11111110;   //*******  
         11'h393: data = 8'b11111110;   //*******
         11'h394: data = 8'b11000110;   //**   **
         11'h395: data = 8'b11000110;   //**   **
         11'h396: data = 8'b11111110;   //*******
         11'h397: data = 8'b11111110;   //*******
         11'h398: data = 8'b00000110;   //     **
         11'h399: data = 8'b00000110;   //     **
         11'h39a: data = 8'b11111110;   //*******
         11'h39b: data = 8'b11111110;   //*******
         11'h39c: data = 8'b00000000;   //
         11'h39d: data = 8'b00000000;   //
         11'h39e: data = 8'b00000000;   //
         11'h39f: data = 8'b00000000;   //
          // code x3a (:)
         11'h3a0: data = 8'b00000000;   //
         11'h3a1: data = 8'b00000000;   //
         11'h3a2: data = 8'b00000000;   //
         11'h3a3: data = 8'b00000000;   //
         11'h3a4: data = 8'b00011000;   //   **
         11'h3a5: data = 8'b00011000;   //   **
         11'h3a6: data = 8'b00000000;   //
         11'h3a7: data = 8'b00000000;   //
         11'h3a8: data = 8'b00011000;   //   **
         11'h3a9: data = 8'b00011000;   //   **
         11'h3aa: data = 8'b00000000;   //   
         11'h3ab: data = 8'b00000000;   //   
         11'h3ac: data = 8'b00000000;   //
         11'h3ad: data = 8'b00000000;   //
         11'h3ae: data = 8'b00000000;   //
         11'h3af: data = 8'b00000000;   //
         // **** MAKE SHIFT ASCII FOR CLOCK / CALENDAR      
         // code x40 (A)
         11'h400: data = 8'b00000000;   //
         11'h401: data = 8'b00000000;   //
         11'h402: data = 8'b00010000;   //   *
         11'h403: data = 8'b00111000;   //  ***
         11'h404: data = 8'b01101100;   // ** **   
         11'h405: data = 8'b11000110;   //**   **   
         11'h406: data = 8'b11000110;   //**   **
         11'h407: data = 8'b11111110;   //*******
         11'h408: data = 8'b11111110;   //*******
         11'h409: data = 8'b11000110;   //**   **
         11'h40a: data = 8'b11000110;   //**   **
         11'h40b: data = 8'b11000110;   //**   **
         11'h40c: data = 8'b00000000;   //
         11'h40d: data = 8'b00000000;   //
         11'h40e: data = 8'b00000000;   //
         11'h40f: data = 8'b00000000;   //
         // code x41 (P)
         11'h410: data = 8'b00000000;   //
         11'h411: data = 8'b00000000;   //
         11'h412: data = 8'b11111100;   //******
         11'h413: data = 8'b11111110;   //*******
         11'h414: data = 8'b11000110;   //**   **
         11'h415: data = 8'b11000110;   //**   **
         11'h416: data = 8'b11111110;   //*******
         11'h417: data = 8'b11111100;   //****** 
         11'h418: data = 8'b11000000;   //**   
         11'h419: data = 8'b11000000;   //**   
         11'h41a: data = 8'b11000000;   //**
         11'h41b: data = 8'b11000000;   //**
         11'h41c: data = 8'b00000000;   //
         11'h41d: data = 8'b00000000;   //
         11'h41e: data = 8'b00000000;   //
         11'h41f: data = 8'b00000000;   //
         // code x4d (M)
         11'h4d0: data = 8'b00000000;   //
         11'h4d1: data = 8'b00000000;   //
         11'h4d2: data = 8'b11000110;   //**   **
         11'h4d3: data = 8'b11000110;   //**   **
         11'h4d4: data = 8'b11101110;   //*** ***
         11'h4d5: data = 8'b11111110;   //*******
         11'h4d6: data = 8'b11010110;   //** * **
         11'h4d7: data = 8'b11000110;   //**   **
         11'h4d8: data = 8'b11000110;   //**   **
         11'h4d9: data = 8'b11000110;   //**   **
         11'h4da: data = 8'b11000110;   //**   **
         11'h4db: data = 8'b11000110;   //**   **
         11'h4dc: data = 8'b00000000;   //
         11'h4dd: data = 8'b00000000;   //
         11'h4de: data = 8'b00000000;   //
         11'h4df: data = 8'b00000000;   //
         
            // code x51 (S)
         11'h510: data = 8'b00000000;   //
         11'h511: data = 8'b00000000;   //
         11'h512: data = 8'b11111110;   //*******
         11'h513: data = 8'b11111110;   //*******   
         11'h514: data = 8'b11000000;   //**   
         11'h515: data = 8'b11000000;   //**
         11'h516: data = 8'b11111110;   //*******
         11'h517: data = 8'b11111110;   //*******
         11'h518: data = 8'b00000110;   //     **
         11'h519: data = 8'b00000110;   //     **
         11'h51a: data = 8'b11111110;   //*******
         11'h51b: data = 8'b11111110;   //*******
         11'h51c: data = 8'b00000000;   //
         11'h51d: data = 8'b00000000;   //
         11'h51e: data = 8'b00000000;   //
         11'h51f: data = 8'b00000000;   //
         
         
            // code x52 (T)
         11'h520: data = 8'b00000000;   //
         11'h521: data = 8'b00000000;   //
         11'h522: data = 8'b11111110;   //******
         11'h523: data = 8'b11111110;   //******   
         11'h524: data = 8'b00011000;   //  **   
         11'h525: data = 8'b00011000;   //  **
         11'h526: data = 8'b00011000;   //  **
         11'h527: data = 8'b00011000;   //  **
         11'h528: data = 8'b00011000;   //  **
         11'h529: data = 8'b00011000;   //  **
         11'h52a: data = 8'b00011000;   //  **
         11'h52b: data = 8'b00011000;   //  **
         11'h52c: data = 8'b00000000;   //
         11'h52d: data = 8'b00000000;   //
         11'h52e: data = 8'b00000000;   //
         11'h52f: data = 8'b00000000;   //
         
          default: data = 8'b00000000;    // default
      endcase
   
endmodule